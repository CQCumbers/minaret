`include "defines.sv"
`include "mfi_testbench.sv"
`include "mfi_pc_fwd_check.sv"
