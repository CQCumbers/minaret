`define MINA_FORMAL
`define MINA_FORMAL_CHECKER mfi_inst_check
`define MINA_FORMAL_RESET_CYCLES 1
`define MINA_FORMAL_CHECK_CYCLE 20
`define MINA_FORMAL_INST_MODEL mfi_inst_add
`define DEBUGNETS
`include "mfi_macros.vh"

