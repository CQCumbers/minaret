`include "defines.sv"
`include "mfi_testbench.sv"
`include "mfi_inst_check.sv"
`include "inst_sub.v"
