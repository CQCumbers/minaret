`define MINA_FORMAL
`define MINA_FORMAL_CHECKER mfi_pc_fwd_check
`define MINA_FORMAL_RESET_CYCLES 10
`define MINA_FORMAL_CHECK_CYCLE 30
`define DEBUGNETS
`include "mfi_macros.vh"

